bind z2_2 z2_2_checker c0(.clk(clk), .rst(rst), .a(a), .b(b), .c(c), .d(d), .e(e), .f(f), .o1(o1), .o2(o2));
