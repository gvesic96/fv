bind z3_all z3_all_checker c0(.clk(clk), 
				.rst(rst), 
				//zadatak1:
				.RT1(RT1),
   				.RDY1(RDY1),
    				.START1(START1),
				.ENDD1(ENDD1),
				//zadatak2:	
				.ER2(ER2),
				//zadatak3:	
				.ER3(ER3),	
				.RDY3(RDY3),
				//zadatak4:
				.RDY4(RDY4),
				.START4(START4),
				//zadatak5:
				.ENDD5(ENDD5),
				.STOP5(STOP5),
				.ER5(ER5),
				.RDY5(RDY5),
				.START5(START5),
				//zadatak6:
				.ENDD6(ENDD6),
				.STOP6(STOP6),
				.ER6(ER6),
				.RDY6(RDY6),
				//zadatak7:
				.ENDD7(ENDD7),
				.START7(START7),
				.STATUS_VALID7(STATUS_VALID7),
				.INSTARTSV7(INSTARTSV7),
				//zadatak8:
				.RT8(RT8),
				.ENABLE8(ENABLE8),
				//zadatak9:
				.RDY9(RDY9),
				.START9(START9),
				.INTERUPT9(INTERUPT9),
				//zadatak10:
				.ACK10(ACK10),
				.REQ10(REQ10));
